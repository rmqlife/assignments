----------------------------------------------------------------------------------
-- Company: 
-- Engineer: 
-- 
-- Create Date:    12:06:04 11/10/2012 
-- Design Name: 
-- Module Name:    instruction_ram - Behavioral 
-- Project Name: 
-- Target Devices: 
-- Tool versions: 
-- Description: 
--
-- Dependencies: 
--
-- Revision: 
-- Revision 0.01 - File Created
-- Additional Comments: 
--
----------------------------------------------------------------------------------
library IEEE;
use IEEE.STD_LOGIC_1164.ALL;

-- Uncomment the following library declaration if using
-- arithmetic functions with Signed or Unsigned values
--use IEEE.NUMERIC_STD.ALL;

-- Uncomment the following library declaration if instantiating
-- any Xilinx primitives in this code.
--library UNISIM;
--use UNISIM.VComponents.all;

entity instruction_ram is
    Port ( pc_in : in  STD_LOGIC_VECTOR (15 downto 0);
           instruction_out : out  STD_LOGIC_VECTOR (15 downto 0);
			  clk : in  STD_LOGIC;
           en : in  STD_LOGIC);
end instruction_ram;

architecture Behavioral of instruction_ram is

begin

end Behavioral;

